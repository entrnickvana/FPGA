`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:33:02 08/26/2017 
// Design Name: 
// Module Name:    led_Mod 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module led_Mod(
	input clock,
	output pins
    );

	always @(posedge clk or posedge rst) 
	begin
		if (rst) 
		begin
			// reset
			
		end
		else if () 
		begin
			
		end
	end


endmodule
